library verilog;
use verilog.vl_types.all;
entity Exercise1Question1 is
    port(
        Y3              : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        Y2              : out    vl_logic;
        Y1              : out    vl_logic;
        Y0              : out    vl_logic
    );
end Exercise1Question1;

library verilog;
use verilog.vl_types.all;
entity Question1_vlg_vec_tst is
end Question1_vlg_vec_tst;

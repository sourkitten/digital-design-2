library verilog;
use verilog.vl_types.all;
entity Exercise1Question1_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Exercise1Question1_vlg_sample_tst;

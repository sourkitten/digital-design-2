library verilog;
use verilog.vl_types.all;
entity MUX16_1_vlg_vec_tst is
end MUX16_1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Question6_vlg_vec_tst is
end Question6_vlg_vec_tst;

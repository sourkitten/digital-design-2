library verilog;
use verilog.vl_types.all;
entity Adder8_vlg_vec_tst is
end Adder8_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Reg8_vlg_vec_tst is
end Reg8_vlg_vec_tst;

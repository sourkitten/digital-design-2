library verilog;
use verilog.vl_types.all;
entity Question4_vlg_vec_tst is
end Question4_vlg_vec_tst;

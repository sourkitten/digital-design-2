library verilog;
use verilog.vl_types.all;
entity Exercise1Question1_vlg_vec_tst is
end Exercise1Question1_vlg_vec_tst;

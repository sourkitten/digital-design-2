library verilog;
use verilog.vl_types.all;
entity Question5_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Question5_vlg_check_tst;

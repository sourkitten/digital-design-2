library verilog;
use verilog.vl_types.all;
entity MUX4_1_vlg_vec_tst is
end MUX4_1_vlg_vec_tst;

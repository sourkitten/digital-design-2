library verilog;
use verilog.vl_types.all;
entity Reg_vlg_vec_tst is
end Reg_vlg_vec_tst;

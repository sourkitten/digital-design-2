library verilog;
use verilog.vl_types.all;
entity Question6_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Question6_vlg_check_tst;

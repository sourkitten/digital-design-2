library verilog;
use verilog.vl_types.all;
entity Exercise1Question3 is
    port(
        F1              : out    vl_logic;
        I2              : in     vl_logic;
        I1              : in     vl_logic;
        I0              : in     vl_logic;
        F0              : out    vl_logic
    );
end Exercise1Question3;

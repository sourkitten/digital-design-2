library verilog;
use verilog.vl_types.all;
entity o8bit_rshifter_loader_vlg_vec_tst is
end o8bit_rshifter_loader_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Question2_vlg_vec_tst is
end Question2_vlg_vec_tst;

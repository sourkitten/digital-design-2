library verilog;
use verilog.vl_types.all;
entity Question5_vlg_vec_tst is
end Question5_vlg_vec_tst;

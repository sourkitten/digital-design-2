library verilog;
use verilog.vl_types.all;
entity Question7_vlg_vec_tst is
end Question7_vlg_vec_tst;
